`ifndef __STATES_VH__

`define __STATES_VH__

`define IDLE 0
`define RUNNING 1
`define SENDING 2
`define PROCESSING_FEW_SHOT 3

`define NUMBER_OF_STATES 4

`endif
